-- FIR filter coefficients
--
-- FI - UAQ
--
-- Electronica Avanzada III
--
-- Rene Romero Troncoso
--

library IEEE;
use IEEE.std_logic_1164.all;

entity ROM is
   port(
      I : in  std_logic_vector(7 downto 0);
      A : out std_logic_vector(23 downto 0)
      );
   end ROM;

architecture LUTable of ROM is
begin
   process(I)
   begin
      case I is
         -- Coefficient format 2.22
         when "00000000" => A <= "000000000011000001100010"; -- Index 0   Coefficient 0.00295305
         when "00000001" => A <= "000000000010111101100101"; -- Index 1   Coefficient 0.00289273
         when "00000010" => A <= "000000000010110001010011"; -- Index 2   Coefficient 0.00270534
         when "00000011" => A <= "000000000010011011011101"; -- Index 3   Coefficient 0.00237203
         when "00000100" => A <= "000000000001111010011100"; -- Index 4   Coefficient 0.00186825
         when "00000101" => A <= "000000000001001100101001"; -- Index 5   Coefficient 0.00116944
         when "00000110" => A <= "000000000000010001000100"; -- Index 6   Coefficient 0.00026035
         when "00000111" => A <= "111111111111000111111001"; -- Index 7   Coefficient -0.00085616
         when "00001000" => A <= "111111111101110010111110"; -- Index 8   Coefficient -0.00215197
         when "00001001" => A <= "111111111100010110001011"; -- Index 9   Coefficient -0.00356793
         when "00001010" => A <= "111111111010110111011100"; -- Index 10   Coefficient -0.00501347
         when "00001011" => A <= "111111111001011110100011"; -- Index 11   Coefficient -0.00636983
         when "00001100" => A <= "111111111000010100101011"; -- Index 12   Coefficient -0.00749707
         when "00001101" => A <= "111111110111100011100111"; -- Index 13   Coefficient -0.00824571
         when "00001110" => A <= "111111110111010100110010"; -- Index 14   Coefficient -0.00847197
         when "00001111" => A <= "111111110111110000001100"; -- Index 15   Coefficient -0.00805378
         when "00010000" => A <= "111111111000111011010001"; -- Index 16   Coefficient -0.00690818
         when "00010001" => A <= "111111111010110111111101"; -- Index 17   Coefficient -0.00500560
         when "00010010" => A <= "111111111101100011111101"; -- Index 18   Coefficient -0.00238109
         when "00010011" => A <= "000000000000111000010100"; -- Index 19   Coefficient 0.00085926
         when "00010100" => A <= "000000000100101001100000"; -- Index 20   Coefficient 0.00453949
         when "00010101" => A <= "000000001000100111110111"; -- Index 21   Coefficient 0.00842071
         when "00010110" => A <= "000000001100100000100010"; -- Index 22   Coefficient 0.01221514
         when "00010111" => A <= "000000001111111110111000"; -- Index 23   Coefficient 0.01560783
         when "00011000" => A <= "000000010010101110000010"; -- Index 24   Coefficient 0.01828051
         when "00011001" => A <= "000000010100011010110011"; -- Index 25   Coefficient 0.01994014
         when "00011010" => A <= "000000010100110101011101"; -- Index 26   Coefficient 0.02034688
         when "00011011" => A <= "000000010011110011011100"; -- Index 27   Coefficient 0.01933956
         when "00011100" => A <= "000000010001010000101101"; -- Index 28   Coefficient 0.01685643
         when "00011101" => A <= "000000001101010000100101"; -- Index 29   Coefficient 0.01294827
         when "00011110" => A <= "000000000111111110001001"; -- Index 30   Coefficient 0.00778413
         when "00011111" => A <= "000000000001101011110011"; -- Index 31   Coefficient 0.00164485
         when "00100000" => A <= "111111111010110010010011"; -- Index 32   Coefficient -0.00509191
         when "00100001" => A <= "111111110011101111001101"; -- Index 33   Coefficient -0.01197505
         when "00100010" => A <= "111111101101000010101110"; -- Index 34   Coefficient -0.01851320
         when "00100011" => A <= "111111100111001101010100"; -- Index 35   Coefficient -0.02421093
         when "00100100" => A <= "111111100010101101000101"; -- Index 36   Coefficient -0.02860904
         when "00100101" => A <= "111111011111111011010100"; -- Index 37   Coefficient -0.03132153
         when "00100110" => A <= "111111011111001010001111"; -- Index 38   Coefficient -0.03207040
         when "00100111" => A <= "111111100000100011010010"; -- Index 39   Coefficient -0.03071165
         when "00101000" => A <= "111111100100000110000001"; -- Index 40   Coefficient -0.02725196
         when "00101001" => A <= "111111101001100111110000"; -- Index 41   Coefficient -0.02185440
         when "00101010" => A <= "111111110000110100001001"; -- Index 42   Coefficient -0.01482940
         when "00101011" => A <= "111111111001001110010110"; -- Index 43   Coefficient -0.00661707
         when "00101100" => A <= "000000000010010011000100"; -- Index 44   Coefficient 0.00224400
         when "00101101" => A <= "000000001011011011000100"; -- Index 45   Coefficient 0.01115513
         when "00101110" => A <= "000000010011111110000110"; -- Index 46   Coefficient 0.01950216
         when "00101111" => A <= "000000011011010101111011"; -- Index 47   Coefficient 0.02670169
         when "00110000" => A <= "111111100100000110000001"; -- Index 40   Coefficient -0.02725196
         when "00110001" => A <= "000000100100100110000111"; -- Index 49   Coefficient 0.03573775
         when "00110010" => A <= "000000100101110100010001"; -- Index 50   Coefficient 0.03693032
         when "00110011" => A <= "000000100100100110000111"; -- Index 51   Coefficient 0.03573775
         when "00110100" => A <= "000000100001000001001101"; -- Index 52   Coefficient 0.03224492
         when "00110101" => A <= "000000011011010101111011"; -- Index 53   Coefficient 0.02670169
         when "00110110" => A <= "000000010011111110000110"; -- Index 54   Coefficient 0.01950216
         when "00110111" => A <= "000000001011011011000100"; -- Index 55   Coefficient 0.01115513
         when "00111000" => A <= "000000000010010011000100"; -- Index 56   Coefficient 0.00224400
         when "00111001" => A <= "111111111001001110010110"; -- Index 57   Coefficient -0.00661707
         when "00111010" => A <= "111111110000110100001001"; -- Index 58   Coefficient -0.01482940
         when "00111011" => A <= "111111101001100111110000"; -- Index 59   Coefficient -0.02185440
         when "00111100" => A <= "111111100100000110000001"; -- Index 60   Coefficient -0.02725196
         when "00111101" => A <= "111111100000100011010010"; -- Index 61   Coefficient -0.03071165
         when "00111110" => A <= "111111011111001010001111"; -- Index 62   Coefficient -0.03207040
         when "00111111" => A <= "111111011111111011010100"; -- Index 63   Coefficient -0.03132153
         when "01000000" => A <= "111111100010101101000101"; -- Index 64   Coefficient -0.02860904
         when "01000001" => A <= "000000011011010101111011"; -- Index 53   Coefficient 0.02670169
         when "01000010" => A <= "111111101101000010101110"; -- Index 66   Coefficient -0.01851320
         when "01000011" => A <= "111111110011101111001101"; -- Index 67   Coefficient -0.01197505
         when "01000100" => A <= "111111111010110010010011"; -- Index 68   Coefficient -0.00509191
         when "01000101" => A <= "000000000001101011110011"; -- Index 69   Coefficient 0.00164485
         when "01000110" => A <= "000000000111111110001001"; -- Index 70   Coefficient 0.00778413
         when "01000111" => A <= "000000001101010000100101"; -- Index 71   Coefficient 0.01294827
         when "01001000" => A <= "000000010001010000101101"; -- Index 72   Coefficient 0.01685643
         when "01001001" => A <= "000000010011110011011100"; -- Index 73   Coefficient 0.01933956
         when "01001010" => A <= "000000010100110101011101"; -- Index 74   Coefficient 0.02034688
         when "01001011" => A <= "000000010100011010110011"; -- Index 75   Coefficient 0.01994014
         when "01001100" => A <= "000000010010101110000010"; -- Index 76   Coefficient 0.01828051
         when "01001101" => A <= "000000001111111110111000"; -- Index 77   Coefficient 0.01560783
         when "01001110" => A <= "000000001100100000100010"; -- Index 78   Coefficient 0.01221514
         when "01001111" => A <= "000000001000100111110111"; -- Index 79   Coefficient 0.00842071
         when "01010000" => A <= "000000000100101001100000"; -- Index 80   Coefficient 0.00453949
         when "01010001" => A <= "000000000000111000010100"; -- Index 81   Coefficient 0.00085926
         when "01010010" => A <= "111111111101100011111101"; -- Index 82   Coefficient -0.00238109
         when "01010011" => A <= "111111111010110111111101"; -- Index 83   Coefficient -0.00500560
         when "01010100" => A <= "111111111000111011010001"; -- Index 84   Coefficient -0.00690818
         when "01010101" => A <= "111111110111110000001100"; -- Index 85   Coefficient -0.00805378
         when "01010110" => A <= "111111110111010100110010"; -- Index 86   Coefficient -0.00847197
         when "01010111" => A <= "111111110111100011100111"; -- Index 87   Coefficient -0.00824571
         when "01011000" => A <= "111111111000010100101011"; -- Index 88   Coefficient -0.00749707
         when "01011001" => A <= "111111111001011110100011"; -- Index 89   Coefficient -0.00636983
         when "01011010" => A <= "111111111010110111011100"; -- Index 90   Coefficient -0.00501347
         when "01011011" => A <= "111111111100010110001011"; -- Index 91   Coefficient -0.00356793
         when "01011100" => A <= "111111111101110010111110"; -- Index 92   Coefficient -0.00215197
         when "01011101" => A <= "111111111111000111111001"; -- Index 93   Coefficient -0.00085616
         when "01011110" => A <= "000000000000010001000100"; -- Index 94   Coefficient 0.00026035
         when "01011111" => A <= "000000000001001100101001"; -- Index 95   Coefficient 0.00116944
         when "01100000" => A <= "000000000001111010011100"; -- Index 96   Coefficient 0.00186825
         when "01100001" => A <= "000000000010011011011101"; -- Index 97   Coefficient 0.00237203
         when "01100010" => A <= "000000000010110001010011"; -- Index 98   Coefficient 0.00270534
         when "01100011" => A <= "000000000010111101100101"; -- Index 99   Coefficient 0.00289273
         when "01100100" => A <= "000000000011000001100010"; -- Index 100   Coefficient 0.00295305
         when others => A <= "000000000000000000000000"; -- Irrelevant indexes
      end case;
   end process;
end LUTable;
